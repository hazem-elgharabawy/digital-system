module edge_bit_counter (
    input counter_enable,
    output edge_count,
    output bit_count
);
    
endmodule