module TOP (
    input           clk,
    input           rst,
    input           PAR_TYP,
    input           PAR_EN,
    input           Prescale,
    input           RX_IN,
    output [10:0]   P_DATA,
    output          data_valid
);
    






    
endmodule