module data_sampling (
    input RX_IN,
    input Prescale,
    input data_sample_en,
    input edge_count,
    output sampled_bit,
);
    
endmodule