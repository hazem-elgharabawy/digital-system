module stop_check (
    input stop_check_en,
    input sampled_bit,
    output stop_err
);
    
endmodule