module parity_check (
    input PAR_TYP,
    input parity_check_en,
    input sampled_bit,
    output par_err
);
    
endmodule