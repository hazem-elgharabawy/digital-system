module start_check (
    input start_check_en,
    input sampled_bit,
    output start_glitch
);
    
endmodule