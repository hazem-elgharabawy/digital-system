module deserializer (
    input sampled_bit,
    input deser_en,
    output P_DATA
);
    
endmodule