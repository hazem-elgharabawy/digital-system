module FSM (
    input PAR_EN,
    input RX_IN,
    input edge_count,
    input bit_count,
    input stop_error
    input start_glitch,
    input par_error,
    output dat_sample_en,
    output counter_enable,
    output deser_en,
    output data_valid,
    output stop_check_en,
    output start_check_en,
    output par_check_en
);


    
endmodule